package counter_pkg;

import uvm_pkg::*;
`include"uvm_macros.svh"

`include "seq_item.sv"
`include "seq.sv"
`include "seqr.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "agent.sv"
`include "environment.sv"
`include "test.sv"

endpackage
